//////////////////////////////////////////////////////////////////////////////////
// Exercise #1 
// Student Name:
// Date: 
//
//  Description: In this exercise, you need to design a logical unit, where the  
//  output acts according to the following truth table:
//
//  a | b | out
// -----------------
//  0 | 0 | func[0]
//  0 | 1 | func [1]
//  1 | 0 | func [2]
//  1 | 1 | func [3]
//
//  inputs:
//           a, b, func[3:0]
//
//  outputs:
//           out
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

module logicalunit(
    input a,
    input b,
    input [3:0] func,
    output out
    );
         
	assign AB = {a, b};  // concatenate a and b bits
	assign out = (AB==2'b00) ? func[0]:
		(AB==2'b01) ? func[1]:
		(AB==2'b10) ? func[2]:
		(AB==2'b11) ? func[3]:
		2'b11;
	

endmodule
